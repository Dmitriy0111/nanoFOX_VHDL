library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.nf_mem_pkg.all;

package nf_program is

    constant program : mem_t(4096*4-1 downto 0)(7 downto 0) :=     (         0 => X"6F",
        1 => X"00",
        2 => X"00",
        3 => X"04",
        4 => X"6F",
        5 => X"00",
        6 => X"80",
        7 => X"11",
        8 => X"6F",
        9 => X"00",
        10 => X"80",
        11 => X"11",
        12 => X"6F",
        13 => X"00",
        14 => X"80",
        15 => X"11",
        16 => X"6F",
        17 => X"00",
        18 => X"80",
        19 => X"11",
        20 => X"6F",
        21 => X"00",
        22 => X"80",
        23 => X"11",
        24 => X"6F",
        25 => X"00",
        26 => X"80",
        27 => X"11",
        28 => X"6F",
        29 => X"00",
        30 => X"80",
        31 => X"11",
        32 => X"6F",
        33 => X"00",
        34 => X"80",
        35 => X"11",
        36 => X"6F",
        37 => X"00",
        38 => X"80",
        39 => X"11",
        40 => X"6F",
        41 => X"00",
        42 => X"80",
        43 => X"11",
        44 => X"6F",
        45 => X"00",
        46 => X"80",
        47 => X"11",
        48 => X"6F",
        49 => X"00",
        50 => X"80",
        51 => X"11",
        52 => X"6F",
        53 => X"00",
        54 => X"80",
        55 => X"11",
        56 => X"6F",
        57 => X"00",
        58 => X"80",
        59 => X"11",
        60 => X"6F",
        61 => X"00",
        62 => X"80",
        63 => X"11",
        64 => X"B7",
        65 => X"00",
        66 => X"00",
        67 => X"00",
        68 => X"37",
        69 => X"01",
        70 => X"00",
        71 => X"00",
        72 => X"B7",
        73 => X"01",
        74 => X"00",
        75 => X"00",
        76 => X"37",
        77 => X"02",
        78 => X"00",
        79 => X"00",
        80 => X"B7",
        81 => X"02",
        82 => X"00",
        83 => X"00",
        84 => X"37",
        85 => X"03",
        86 => X"00",
        87 => X"00",
        88 => X"B7",
        89 => X"03",
        90 => X"00",
        91 => X"00",
        92 => X"37",
        93 => X"04",
        94 => X"00",
        95 => X"00",
        96 => X"B7",
        97 => X"04",
        98 => X"00",
        99 => X"00",
        100 => X"37",
        101 => X"05",
        102 => X"00",
        103 => X"00",
        104 => X"B7",
        105 => X"05",
        106 => X"00",
        107 => X"00",
        108 => X"37",
        109 => X"06",
        110 => X"00",
        111 => X"00",
        112 => X"B7",
        113 => X"06",
        114 => X"00",
        115 => X"00",
        116 => X"37",
        117 => X"07",
        118 => X"00",
        119 => X"00",
        120 => X"B7",
        121 => X"07",
        122 => X"00",
        123 => X"00",
        124 => X"37",
        125 => X"08",
        126 => X"00",
        127 => X"00",
        128 => X"B7",
        129 => X"08",
        130 => X"00",
        131 => X"00",
        132 => X"37",
        133 => X"09",
        134 => X"00",
        135 => X"00",
        136 => X"B7",
        137 => X"09",
        138 => X"00",
        139 => X"00",
        140 => X"37",
        141 => X"0A",
        142 => X"00",
        143 => X"00",
        144 => X"B7",
        145 => X"0A",
        146 => X"00",
        147 => X"00",
        148 => X"37",
        149 => X"0B",
        150 => X"00",
        151 => X"00",
        152 => X"B7",
        153 => X"0B",
        154 => X"00",
        155 => X"00",
        156 => X"37",
        157 => X"0C",
        158 => X"00",
        159 => X"00",
        160 => X"B7",
        161 => X"0C",
        162 => X"00",
        163 => X"00",
        164 => X"37",
        165 => X"0D",
        166 => X"00",
        167 => X"00",
        168 => X"B7",
        169 => X"0D",
        170 => X"00",
        171 => X"00",
        172 => X"37",
        173 => X"0E",
        174 => X"00",
        175 => X"00",
        176 => X"B7",
        177 => X"0E",
        178 => X"00",
        179 => X"00",
        180 => X"37",
        181 => X"0F",
        182 => X"00",
        183 => X"00",
        184 => X"B7",
        185 => X"0F",
        186 => X"00",
        187 => X"00",
        188 => X"37",
        189 => X"11",
        190 => X"00",
        191 => X"00",
        192 => X"13",
        193 => X"01",
        194 => X"01",
        195 => X"00",
        196 => X"6F",
        197 => X"00",
        198 => X"40",
        199 => X"00",
        200 => X"B7",
        201 => X"07",
        202 => X"03",
        203 => X"00",
        204 => X"13",
        205 => X"07",
        206 => X"20",
        207 => X"1B",
        208 => X"23",
        209 => X"A6",
        210 => X"E7",
        211 => X"00",
        212 => X"13",
        213 => X"07",
        214 => X"40",
        215 => X"00",
        216 => X"23",
        217 => X"A0",
        218 => X"E7",
        219 => X"00",
        220 => X"13",
        221 => X"06",
        222 => X"80",
        223 => X"15",
        224 => X"13",
        225 => X"05",
        226 => X"86",
        227 => X"03",
        228 => X"37",
        229 => X"07",
        230 => X"03",
        231 => X"00",
        232 => X"93",
        233 => X"06",
        234 => X"50",
        235 => X"00",
        236 => X"93",
        237 => X"85",
        238 => X"06",
        239 => X"00",
        240 => X"83",
        241 => X"27",
        242 => X"06",
        243 => X"00",
        244 => X"23",
        245 => X"22",
        246 => X"F7",
        247 => X"00",
        248 => X"23",
        249 => X"20",
        250 => X"B7",
        251 => X"00",
        252 => X"83",
        253 => X"27",
        254 => X"07",
        255 => X"00",
        256 => X"E3",
        257 => X"8E",
        258 => X"D7",
        259 => X"FE",
        260 => X"13",
        261 => X"06",
        262 => X"46",
        263 => X"00",
        264 => X"E3",
        265 => X"14",
        266 => X"A6",
        267 => X"FE",
        268 => X"B7",
        269 => X"07",
        270 => X"01",
        271 => X"00",
        272 => X"13",
        273 => X"07",
        274 => X"50",
        275 => X"05",
        276 => X"23",
        277 => X"A2",
        278 => X"E7",
        279 => X"00",
        280 => X"6F",
        281 => X"00",
        282 => X"00",
        283 => X"00",
        284 => X"6F",
        285 => X"00",
        286 => X"00",
        287 => X"00",
        288 => X"6F",
        289 => X"00",
        290 => X"00",
        291 => X"00",
        292 => X"6F",
        293 => X"00",
        294 => X"00",
        295 => X"00",
        296 => X"6F",
        297 => X"00",
        298 => X"00",
        299 => X"00",
        300 => X"6F",
        301 => X"00",
        302 => X"00",
        303 => X"00",
        304 => X"6F",
        305 => X"00",
        306 => X"00",
        307 => X"00",
        308 => X"6F",
        309 => X"00",
        310 => X"00",
        311 => X"00",
        312 => X"6F",
        313 => X"00",
        314 => X"00",
        315 => X"00",
        316 => X"6F",
        317 => X"00",
        318 => X"00",
        319 => X"00",
        320 => X"6F",
        321 => X"00",
        322 => X"00",
        323 => X"00",
        324 => X"6F",
        325 => X"00",
        326 => X"00",
        327 => X"00",
        328 => X"6F",
        329 => X"00",
        330 => X"00",
        331 => X"00",
        332 => X"6F",
        333 => X"00",
        334 => X"00",
        335 => X"00",
        336 => X"6F",
        337 => X"00",
        338 => X"00",
        339 => X"00",
        340 => X"6F",
        341 => X"00",
        342 => X"00",
        343 => X"00",
        344 => X"48",
        345 => X"00",
        346 => X"00",
        347 => X"00",
        348 => X"65",
        349 => X"00",
        350 => X"00",
        351 => X"00",
        352 => X"6C",
        353 => X"00",
        354 => X"00",
        355 => X"00",
        356 => X"6C",
        357 => X"00",
        358 => X"00",
        359 => X"00",
        360 => X"6F",
        361 => X"00",
        362 => X"00",
        363 => X"00",
        364 => X"20",
        365 => X"00",
        366 => X"00",
        367 => X"00",
        368 => X"57",
        369 => X"00",
        370 => X"00",
        371 => X"00",
        372 => X"6F",
        373 => X"00",
        374 => X"00",
        375 => X"00",
        376 => X"72",
        377 => X"00",
        378 => X"00",
        379 => X"00",
        380 => X"6C",
        381 => X"00",
        382 => X"00",
        383 => X"00",
        384 => X"64",
        385 => X"00",
        386 => X"00",
        387 => X"00",
        388 => X"21",
        389 => X"00",
        390 => X"00",
        391 => X"00",
        392 => X"0A",
        393 => X"00",
        394 => X"00",
        395 => X"00",
        396 => X"0D",
        397 => X"00",
        398 => X"00",
        399 => X"00",
        others => X"XX"
    );

end package nf_program;
