library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.nf_mem_pkg.all;

package nf_program is

    constant program : mem_t(4096*4-1 downto 0)(7 downto 0) :=     (         0 => X"6F",
        1 => X"00",
        2 => X"00",
        3 => X"04",
        4 => X"6F",
        5 => X"00",
        6 => X"00",
        7 => X"0F",
        8 => X"6F",
        9 => X"00",
        10 => X"00",
        11 => X"0F",
        12 => X"6F",
        13 => X"00",
        14 => X"00",
        15 => X"0F",
        16 => X"6F",
        17 => X"00",
        18 => X"00",
        19 => X"0F",
        20 => X"6F",
        21 => X"00",
        22 => X"00",
        23 => X"0F",
        24 => X"6F",
        25 => X"00",
        26 => X"00",
        27 => X"0F",
        28 => X"6F",
        29 => X"00",
        30 => X"00",
        31 => X"0F",
        32 => X"6F",
        33 => X"00",
        34 => X"00",
        35 => X"0F",
        36 => X"6F",
        37 => X"00",
        38 => X"00",
        39 => X"0F",
        40 => X"6F",
        41 => X"00",
        42 => X"00",
        43 => X"0F",
        44 => X"6F",
        45 => X"00",
        46 => X"00",
        47 => X"0F",
        48 => X"6F",
        49 => X"00",
        50 => X"00",
        51 => X"0F",
        52 => X"6F",
        53 => X"00",
        54 => X"00",
        55 => X"0F",
        56 => X"6F",
        57 => X"00",
        58 => X"00",
        59 => X"0F",
        60 => X"6F",
        61 => X"00",
        62 => X"00",
        63 => X"0F",
        64 => X"B7",
        65 => X"00",
        66 => X"00",
        67 => X"00",
        68 => X"37",
        69 => X"01",
        70 => X"00",
        71 => X"00",
        72 => X"B7",
        73 => X"01",
        74 => X"00",
        75 => X"00",
        76 => X"37",
        77 => X"02",
        78 => X"00",
        79 => X"00",
        80 => X"B7",
        81 => X"02",
        82 => X"00",
        83 => X"00",
        84 => X"37",
        85 => X"03",
        86 => X"00",
        87 => X"00",
        88 => X"B7",
        89 => X"03",
        90 => X"00",
        91 => X"00",
        92 => X"37",
        93 => X"04",
        94 => X"00",
        95 => X"00",
        96 => X"B7",
        97 => X"04",
        98 => X"00",
        99 => X"00",
        100 => X"37",
        101 => X"05",
        102 => X"00",
        103 => X"00",
        104 => X"B7",
        105 => X"05",
        106 => X"00",
        107 => X"00",
        108 => X"37",
        109 => X"06",
        110 => X"00",
        111 => X"00",
        112 => X"B7",
        113 => X"06",
        114 => X"00",
        115 => X"00",
        116 => X"37",
        117 => X"07",
        118 => X"00",
        119 => X"00",
        120 => X"B7",
        121 => X"07",
        122 => X"00",
        123 => X"00",
        124 => X"37",
        125 => X"08",
        126 => X"00",
        127 => X"00",
        128 => X"B7",
        129 => X"08",
        130 => X"00",
        131 => X"00",
        132 => X"37",
        133 => X"09",
        134 => X"00",
        135 => X"00",
        136 => X"B7",
        137 => X"09",
        138 => X"00",
        139 => X"00",
        140 => X"37",
        141 => X"0A",
        142 => X"00",
        143 => X"00",
        144 => X"B7",
        145 => X"0A",
        146 => X"00",
        147 => X"00",
        148 => X"37",
        149 => X"0B",
        150 => X"00",
        151 => X"00",
        152 => X"B7",
        153 => X"0B",
        154 => X"00",
        155 => X"00",
        156 => X"37",
        157 => X"0C",
        158 => X"00",
        159 => X"00",
        160 => X"B7",
        161 => X"0C",
        162 => X"00",
        163 => X"00",
        164 => X"37",
        165 => X"0D",
        166 => X"00",
        167 => X"00",
        168 => X"B7",
        169 => X"0D",
        170 => X"00",
        171 => X"00",
        172 => X"37",
        173 => X"0E",
        174 => X"00",
        175 => X"00",
        176 => X"B7",
        177 => X"0E",
        178 => X"00",
        179 => X"00",
        180 => X"37",
        181 => X"0F",
        182 => X"00",
        183 => X"00",
        184 => X"B7",
        185 => X"0F",
        186 => X"00",
        187 => X"00",
        188 => X"37",
        189 => X"11",
        190 => X"00",
        191 => X"00",
        192 => X"13",
        193 => X"01",
        194 => X"01",
        195 => X"00",
        196 => X"6F",
        197 => X"00",
        198 => X"40",
        199 => X"00",
        200 => X"13",
        201 => X"01",
        202 => X"01",
        203 => X"FF",
        204 => X"23",
        205 => X"26",
        206 => X"01",
        207 => X"00",
        208 => X"13",
        209 => X"07",
        210 => X"10",
        211 => X"00",
        212 => X"93",
        213 => X"07",
        214 => X"10",
        215 => X"00",
        216 => X"B3",
        217 => X"87",
        218 => X"E7",
        219 => X"00",
        220 => X"93",
        221 => X"87",
        222 => X"17",
        223 => X"00",
        224 => X"23",
        225 => X"26",
        226 => X"F1",
        227 => X"00",
        228 => X"83",
        229 => X"26",
        230 => X"C1",
        231 => X"00",
        232 => X"93",
        233 => X"07",
        234 => X"07",
        235 => X"00",
        236 => X"13",
        237 => X"87",
        238 => X"06",
        239 => X"00",
        240 => X"6F",
        241 => X"F0",
        242 => X"9F",
        243 => X"FE",
        244 => X"6F",
        245 => X"00",
        246 => X"00",
        247 => X"00",
        248 => X"6F",
        249 => X"00",
        250 => X"00",
        251 => X"00",
        252 => X"6F",
        253 => X"00",
        254 => X"00",
        255 => X"00",
        256 => X"6F",
        257 => X"00",
        258 => X"00",
        259 => X"00",
        260 => X"6F",
        261 => X"00",
        262 => X"00",
        263 => X"00",
        264 => X"6F",
        265 => X"00",
        266 => X"00",
        267 => X"00",
        268 => X"6F",
        269 => X"00",
        270 => X"00",
        271 => X"00",
        272 => X"6F",
        273 => X"00",
        274 => X"00",
        275 => X"00",
        276 => X"6F",
        277 => X"00",
        278 => X"00",
        279 => X"00",
        280 => X"6F",
        281 => X"00",
        282 => X"00",
        283 => X"00",
        284 => X"6F",
        285 => X"00",
        286 => X"00",
        287 => X"00",
        288 => X"6F",
        289 => X"00",
        290 => X"00",
        291 => X"00",
        292 => X"6F",
        293 => X"00",
        294 => X"00",
        295 => X"00",
        296 => X"6F",
        297 => X"00",
        298 => X"00",
        299 => X"00",
        300 => X"6F",
        301 => X"00",
        302 => X"00",
        303 => X"00",
        others => X"XX"
    );

end package nf_program;
