library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.nf_mem_pkg.all;

package nf_program is

    constant program : mem_t(4096*4-1 downto 0)(7 downto 0) :=     (         0 => X"6F",
        1 => X"00",
        2 => X"00",
        3 => X"04",
        4 => X"6F",
        5 => X"00",
        6 => X"C0",
        7 => X"13",
        8 => X"6F",
        9 => X"00",
        10 => X"C0",
        11 => X"13",
        12 => X"6F",
        13 => X"00",
        14 => X"C0",
        15 => X"13",
        16 => X"6F",
        17 => X"00",
        18 => X"C0",
        19 => X"13",
        20 => X"6F",
        21 => X"00",
        22 => X"C0",
        23 => X"13",
        24 => X"6F",
        25 => X"00",
        26 => X"C0",
        27 => X"13",
        28 => X"6F",
        29 => X"00",
        30 => X"C0",
        31 => X"13",
        32 => X"6F",
        33 => X"00",
        34 => X"C0",
        35 => X"13",
        36 => X"6F",
        37 => X"00",
        38 => X"C0",
        39 => X"13",
        40 => X"6F",
        41 => X"00",
        42 => X"C0",
        43 => X"13",
        44 => X"6F",
        45 => X"00",
        46 => X"C0",
        47 => X"13",
        48 => X"6F",
        49 => X"00",
        50 => X"C0",
        51 => X"13",
        52 => X"6F",
        53 => X"00",
        54 => X"C0",
        55 => X"13",
        56 => X"6F",
        57 => X"00",
        58 => X"C0",
        59 => X"13",
        60 => X"6F",
        61 => X"00",
        62 => X"C0",
        63 => X"13",
        64 => X"B7",
        65 => X"00",
        66 => X"00",
        67 => X"00",
        68 => X"37",
        69 => X"01",
        70 => X"00",
        71 => X"00",
        72 => X"B7",
        73 => X"01",
        74 => X"00",
        75 => X"00",
        76 => X"37",
        77 => X"02",
        78 => X"00",
        79 => X"00",
        80 => X"B7",
        81 => X"02",
        82 => X"00",
        83 => X"00",
        84 => X"37",
        85 => X"03",
        86 => X"00",
        87 => X"00",
        88 => X"B7",
        89 => X"03",
        90 => X"00",
        91 => X"00",
        92 => X"37",
        93 => X"04",
        94 => X"00",
        95 => X"00",
        96 => X"B7",
        97 => X"04",
        98 => X"00",
        99 => X"00",
        100 => X"37",
        101 => X"05",
        102 => X"00",
        103 => X"00",
        104 => X"B7",
        105 => X"05",
        106 => X"00",
        107 => X"00",
        108 => X"37",
        109 => X"06",
        110 => X"00",
        111 => X"00",
        112 => X"B7",
        113 => X"06",
        114 => X"00",
        115 => X"00",
        116 => X"37",
        117 => X"07",
        118 => X"00",
        119 => X"00",
        120 => X"B7",
        121 => X"07",
        122 => X"00",
        123 => X"00",
        124 => X"37",
        125 => X"08",
        126 => X"00",
        127 => X"00",
        128 => X"B7",
        129 => X"08",
        130 => X"00",
        131 => X"00",
        132 => X"37",
        133 => X"09",
        134 => X"00",
        135 => X"00",
        136 => X"B7",
        137 => X"09",
        138 => X"00",
        139 => X"00",
        140 => X"37",
        141 => X"0A",
        142 => X"00",
        143 => X"00",
        144 => X"B7",
        145 => X"0A",
        146 => X"00",
        147 => X"00",
        148 => X"37",
        149 => X"0B",
        150 => X"00",
        151 => X"00",
        152 => X"B7",
        153 => X"0B",
        154 => X"00",
        155 => X"00",
        156 => X"37",
        157 => X"0C",
        158 => X"00",
        159 => X"00",
        160 => X"B7",
        161 => X"0C",
        162 => X"00",
        163 => X"00",
        164 => X"37",
        165 => X"0D",
        166 => X"00",
        167 => X"00",
        168 => X"B7",
        169 => X"0D",
        170 => X"00",
        171 => X"00",
        172 => X"37",
        173 => X"0E",
        174 => X"00",
        175 => X"00",
        176 => X"B7",
        177 => X"0E",
        178 => X"00",
        179 => X"00",
        180 => X"37",
        181 => X"0F",
        182 => X"00",
        183 => X"00",
        184 => X"B7",
        185 => X"0F",
        186 => X"00",
        187 => X"00",
        188 => X"37",
        189 => X"11",
        190 => X"00",
        191 => X"00",
        192 => X"13",
        193 => X"01",
        194 => X"01",
        195 => X"00",
        196 => X"6F",
        197 => X"00",
        198 => X"80",
        199 => X"02",
        200 => X"23",
        201 => X"2E",
        202 => X"A0",
        203 => X"16",
        204 => X"83",
        205 => X"27",
        206 => X"C0",
        207 => X"17",
        208 => X"63",
        209 => X"8C",
        210 => X"07",
        211 => X"00",
        212 => X"83",
        213 => X"27",
        214 => X"C0",
        215 => X"17",
        216 => X"93",
        217 => X"87",
        218 => X"F7",
        219 => X"FF",
        220 => X"23",
        221 => X"2E",
        222 => X"F0",
        223 => X"16",
        224 => X"83",
        225 => X"27",
        226 => X"C0",
        227 => X"17",
        228 => X"E3",
        229 => X"98",
        230 => X"07",
        231 => X"FE",
        232 => X"67",
        233 => X"80",
        234 => X"00",
        235 => X"00",
        236 => X"13",
        237 => X"01",
        238 => X"01",
        239 => X"FF",
        240 => X"23",
        241 => X"26",
        242 => X"11",
        243 => X"00",
        244 => X"23",
        245 => X"24",
        246 => X"81",
        247 => X"00",
        248 => X"23",
        249 => X"22",
        250 => X"91",
        251 => X"00",
        252 => X"23",
        253 => X"20",
        254 => X"21",
        255 => X"01",
        256 => X"B7",
        257 => X"07",
        258 => X"01",
        259 => X"00",
        260 => X"13",
        261 => X"07",
        262 => X"10",
        263 => X"00",
        264 => X"23",
        265 => X"A2",
        266 => X"E7",
        267 => X"00",
        268 => X"37",
        269 => X"04",
        270 => X"01",
        271 => X"00",
        272 => X"13",
        273 => X"09",
        274 => X"40",
        275 => X"01",
        276 => X"93",
        277 => X"04",
        278 => X"00",
        279 => X"00",
        280 => X"6F",
        281 => X"00",
        282 => X"00",
        283 => X"01",
        284 => X"83",
        285 => X"27",
        286 => X"04",
        287 => X"00",
        288 => X"B3",
        289 => X"07",
        290 => X"F7",
        291 => X"00",
        292 => X"23",
        293 => X"22",
        294 => X"F4",
        295 => X"00",
        296 => X"13",
        297 => X"05",
        298 => X"A0",
        299 => X"00",
        300 => X"EF",
        301 => X"F0",
        302 => X"DF",
        303 => X"F9",
        304 => X"03",
        305 => X"27",
        306 => X"44",
        307 => X"00",
        308 => X"93",
        309 => X"87",
        310 => X"04",
        311 => X"00",
        312 => X"E3",
        313 => X"12",
        314 => X"27",
        315 => X"FF",
        316 => X"6F",
        317 => X"F0",
        318 => X"9F",
        319 => X"FE",
        320 => X"6F",
        321 => X"00",
        322 => X"00",
        323 => X"00",
        324 => X"6F",
        325 => X"00",
        326 => X"00",
        327 => X"00",
        328 => X"6F",
        329 => X"00",
        330 => X"00",
        331 => X"00",
        332 => X"6F",
        333 => X"00",
        334 => X"00",
        335 => X"00",
        336 => X"6F",
        337 => X"00",
        338 => X"00",
        339 => X"00",
        340 => X"6F",
        341 => X"00",
        342 => X"00",
        343 => X"00",
        344 => X"6F",
        345 => X"00",
        346 => X"00",
        347 => X"00",
        348 => X"6F",
        349 => X"00",
        350 => X"00",
        351 => X"00",
        352 => X"6F",
        353 => X"00",
        354 => X"00",
        355 => X"00",
        356 => X"6F",
        357 => X"00",
        358 => X"00",
        359 => X"00",
        360 => X"6F",
        361 => X"00",
        362 => X"00",
        363 => X"00",
        364 => X"6F",
        365 => X"00",
        366 => X"00",
        367 => X"00",
        368 => X"6F",
        369 => X"00",
        370 => X"00",
        371 => X"00",
        372 => X"6F",
        373 => X"00",
        374 => X"00",
        375 => X"00",
        376 => X"6F",
        377 => X"00",
        378 => X"00",
        379 => X"00",
        others => X"XX"
    );

end package nf_program;
