/*
*  File            :   nf_tb.svh
*  Autor           :   Vlasov D.V.
*  Data            :   2018.11.28
*  Language        :   SystemVerilog
*  Description     :   This is testbench header for cpu unit
*  Copyright(c)    :   2018 - 2019 Vlasov D.V.
*/

// enable debug instruction messages
`define debug_lev0  0
// enable term logging
`define log_term    1
// enable txt logging
`define log_txt     1
// enable html logging
`define log_html    0
// enable logging
`define log_en      1
